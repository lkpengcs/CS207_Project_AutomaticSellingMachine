`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 2020/12/22 20:13:56
// Design Name: 
// Module Name: top_design
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 2020/12/19 19:11:03
// Design Name: 
// Module Name: top_design
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module top_design(
//basic
input clk,//clock
input rst,//reset
input [3:0] row_data,//used for matrix keyboard input
output [3:0]col_data,//used for matrix keyboard input
//query state
input shift1,shift2,shift3,shift4,//select goods channel
input inenter_pay,//enter pay state
output beep,//output for buzzer
//paying state
input inmoney1,inmoney2,inmoney3,inmoney4,//four kinds of money
input ins1,ins2,ins3,ins4,//select four items when paying
output [6:0] led_en,//status signal (led) for paying
//manager state
input chd1,chd2,chd3,chd4,//the aisle chosen for replenishment
input csw1,//query the quantity sold
input csw2,//supplement goods
input csw3,//query the total price
input inmanager,//to enter manager state
input in_manager_rst,//reset signal for manager

output reg [7:0] segment_led,//seven segment digital tube
output reg [7:0] seg_en//enable signal for seven segment digital tube

    );
//3 different states    
parameter [1:0] state_st=2'b00,state_query=2'b01,state_pay=2'b10,state_manager=2'b11;
reg [1:0] state;
//3 different clock generated by frequency divider
wire clkout1,clkout2,clkout3;
frequency_divider #(100_000_000)u_divider1(clk,rst,clkout1);
frequency_divider #(100_000)u_divider2(clk,rst,clkout2);
frequency_divider #(200_000_000)u_divider3(clk,rst,clkout3);
//seven segment digital tube and enable signal generated by three separated modules
wire [7:0] segment_led1,segment_led2,segment_led3;
wire [7:0] seg_en1,seg_en2,seg_en3;

wire flag;//whether the payment is successful, 1 for true

reg rst1,rst2;//reset signal for query state and paying state

wire[3:0]key_value;//key value output by matrix keyboard
matrix_input u_matrix_input(clk,rst,row_data,key_value,col_data);

wire enter_pay;//whether to enter payment, 1 for true
debounce u_enter_pay(clk,rst,inenter_pay,enter_pay);

wire manager;//enter manager state signal after debounce
debounce u_manager(clk,rst,inmanager,manager);

wire manager_rst;//reset signal for manager after debounce
debounce u_manager_rst(clk,rst,in_manager_rst,manager_rst);

reg [7:0] in1num1,in1num2,in1num3,in1num4;//the number of items before replenishment
wire [7:0] out1num1,out1num2,out1num3,out1num4;//the number of items after replenishment
reg [7:0] in2num1,in2num2,in2num3,in2num4;//the number of items before pay
wire [7:0] out2num1,out2num2,out2num3,out2num4;//the number of items after pay
wire [7:0] require_money;//money needed during one payment, money earned by one payment
wire[7:0] sellnum1,sellnum2,sellnum3,sellnum4;//The quantity of each item sold each time
reg [7:0] in_S1_sell,in_S2_sell,in_S3_sell,in_S4_sell;//The quantity of each item having been sold
reg [7:0] price_sum;//total sales

//initialization
initial begin
state=state_st;
in1num1=8'd0;
in1num2=8'd0;
in1num3=8'd0;
in1num4=8'd0;
in2num1=8'd0;
in2num2=8'd0;
in2num3=8'd0;
in2num4=8'd0;
rst1=1'b0;
rst2=1'b0;
in_S1_sell=8'd0;
in_S2_sell=8'd0;
in_S3_sell=8'd0;
in_S4_sell=8'd0;
price_sum=8'd0;
end

//instantiate three main modules
query u_module_1(clk,clkout1,clkout2,rst1,enter_pay,shift1,shift2,shift3,shift4,
in1num1,in1num2,in1num3,in1num4,
seg_en1,segment_led1,
beep);

paying u_module_2(clk,clkout1,clkout2,clkout3,rst2,
key_value,
inmoney1,inmoney2,inmoney3,inmoney4,
ins1,ins2,ins3,ins4,
in2num1,in2num2,in2num3,in2num4,
out2num1,out2num2,out2num3,out2num4,
segment_led2,
seg_en2,
led_en,
require_money,sellnum1,sellnum2,sellnum3,sellnum4,flag);

replenishment u_module_3(clk,clkout1,clkout2,
manager_rst,
chd1,chd2,chd3,chd4,
csw1,
csw2,
csw3,
key_value,
seg_en3,
segment_led3,
in_S1_sell,in_S2_sell,in_S3_sell,in_S4_sell,
in1num1,in1num2,in1num3,in1num4,
price_sum,
out1num1,out1num2,out1num3,out1num4
      );

//FSM
always @ (negedge clkout2)
begin
    if(!rst)//initialization
    begin     
        state=state_st;
        segment_led=8'b1111_1111;
        seg_en=8'b1111_1111;
        in1num1=8'd0;
        in1num2=8'd0;
        in1num3=8'd0;
        in1num4=8'd0;
        in2num1=8'd0;
        in2num2=8'd0;
        in2num3=8'd0;
        in2num4=8'd0;        
        rst1=1'b0;
        rst2=1'b0;
        in_S1_sell=8'd0;
        in_S2_sell=8'd0;
        in_S3_sell=8'd0;
        in_S4_sell=8'd0;
        price_sum=8'd0;
    end
    else
    begin
    case(state)
    state_st:
    begin
        in1num1=in1num1;
        in1num2=in1num2;
        in1num3=in1num3;
        in1num4=in1num4;
        in2num1=in2num1;
        in2num2=in2num2;
        in2num3=in2num3;
        in2num4=in2num4; 
        segment_led=segment_led;
        seg_en=seg_en;    
        in_S1_sell=in_S1_sell;
        in_S2_sell=in_S2_sell;
        in_S3_sell=in_S3_sell;
        in_S4_sell=in_S4_sell;   
        price_sum=price_sum;//keep every variable unchanged
        if(manager)//enter manager state
        begin
            rst1=1'b0;
            rst2=1'b0;
            state=state_manager;
        end
        else
        begin
            rst1=1'b1;
            rst2=1'b0;
            state=state_query;        
        end   
    end
    
    state_query:
    begin
        if(manager)//enter manager state
        begin
            rst1=1'b0;
            rst2=1'b0;
            state=state_manager;
        end
        else
        begin    
            segment_led=segment_led1;
            seg_en=seg_en1;  
            if(enter_pay)//enter pay state
            begin
                rst1=1'b0;
                rst2=1'b1;        
                state=state_pay;
            end
            else
            begin
                state=state_query;
            end       
        end     

    end
    
    state_pay:
    begin
        if(manager)//enter manager state
        begin
            rst1=1'b0;
            rst2=1'b0;
            state=state_manager;
        end
        else
        begin
            segment_led=segment_led2;
            seg_en=seg_en2;
            if(flag)//payment is successful, then update related variable     
            begin
            in1num1=out2num1;
            in1num2=out2num2;
            in1num3=out2num3;
            in1num4=out2num4;
            in_S1_sell=in_S1_sell+sellnum1;
            in_S2_sell=in_S2_sell+sellnum2;
            in_S3_sell=in_S3_sell+sellnum3;
            in_S4_sell=in_S4_sell+sellnum4;
            price_sum=price_sum+require_money;            
            in2num1=out2num1;
            in2num2=out2num2;
            in2num3=out2num3;
            in2num4=out2num4;            
            end     
            else
            begin
            in1num1=in1num1;
            in1num2=in1num2;
            in1num3=in1num3;
            in1num4=in1num4;
            in_S1_sell=in_S1_sell;
            in_S2_sell=in_S2_sell;
            in_S3_sell=in_S3_sell;
            in_S4_sell=in_S4_sell;
            price_sum=price_sum;            
            in2num1=in2num1;
            in2num2=in2num2;
            in2num3=in2num3;
            in2num4=in2num4;              
            end
            if(!enter_pay)//enter query state
            begin
                rst1=1'b1;
                rst2=1'b0;        
                state=state_query;
            end
            else
            begin
                state=state_pay;
            end  
        end      
    end
    
    state_manager:
    begin
        segment_led=segment_led3;
        seg_en=seg_en3;
        in2num1=out1num1;//update related variable after replenishment
        in2num2=out1num2;
        in2num3=out1num3;
        in2num4=out1num4;
        in1num1=out1num1;
        in1num2=out1num2;
        in1num3=out1num3;
        in1num4=out1num4; 
        in_S1_sell=in_S1_sell;
        in_S2_sell=in_S2_sell;
        in_S3_sell=in_S3_sell;
        in_S4_sell=in_S4_sell;
        price_sum=price_sum;                
        if(!manager)//enter query state
        begin
            rst1=1'b1;
            rst2=1'b0;
            state=state_query;
        end
        else
        begin 
            state=state_manager;        
        end
    end
    endcase
    end
end
endmodule

